`timescale 1ns/1ps

module instruction_mem #(parameter BRAM_ADDR_WIDTH = 10, BRAM_DATA_WIDTH = 32) (clk, addr, wr_n, rd_n, bram_data_out);

    input clk, wr_n, rd_n;
    input [BRAM_ADDR_WIDTH-1:0] addr;
    output reg [BRAM_DATA_WIDTH-1:0] bram_data_out;

    reg [BRAM_DATA_WIDTH-1:0] mem [(1<<BRAM_ADDR_WIDTH)-1:0];
    integer i;
    initial begin
        $monitor("ins mem[%d] = %d at %d", 0, mem[0], $time);
        $readmemb("instructions.mem", mem);
    end

    always @(posedge clk) begin
        if (rd_n == 1'b1) bram_data_out <= mem[addr];
    end

endmodule